module BinaryBCD (
	input [6:0] binary_in,
	output [7:0] bcd_out
);

always_comb
	case (binary_in)
		7'b0000000: bcd_out<= 8'b00000000;
		7'b0000001: bcd_out<= 8'b00000001;
		7'b0000010: bcd_out<= 8'b00000010;
		7'b0000011: bcd_out<= 8'b00000011;
		7'b0000100: bcd_out<= 8'b00000100;
		7'b0000101: bcd_out<= 8'b00000101;
		7'b0000110: bcd_out<= 8'b00000110;
		7'b0000111: bcd_out<= 8'b00000111;
		7'b0001000: bcd_out<= 8'b00001000;
		7'b0001001: bcd_out<= 8'b00001001;
		7'b0001010: bcd_out<= 8'b00010000;
		7'b0001011: bcd_out<= 8'b00010001;
		7'b0001100: bcd_out<= 8'b00010010;
		7'b0001101: bcd_out<= 8'b00010011;
		7'b0001110: bcd_out<= 8'b00010100;
		7'b0001111: bcd_out<= 8'b00010101;
		7'b0010000: bcd_out<= 8'b00010110;
		7'b0010001: bcd_out<= 8'b00010111;
		7'b0010010: bcd_out<= 8'b00011000;
		7'b0010011: bcd_out<= 8'b00011001;
		7'b0010100: bcd_out<= 8'b00100000;
		7'b0010101: bcd_out<= 8'b00100001;
		7'b0010110: bcd_out<= 8'b00100010;
		7'b0010111: bcd_out<= 8'b00100011;
		7'b0011000: bcd_out<= 8'b00100100;
		7'b0011001: bcd_out<= 8'b00100101;
		7'b0011010: bcd_out<= 8'b00100110;
		7'b0011011: bcd_out<= 8'b00100111;
		7'b0011100: bcd_out<= 8'b00101000;
		7'b0011101: bcd_out<= 8'b00101001;
		7'b0011110: bcd_out<= 8'b00110000;
		7'b0011111: bcd_out<= 8'b00110001;
		7'b0100000: bcd_out<= 8'b00110010;
		7'b0100001: bcd_out<= 8'b00110011;
		7'b0100010: bcd_out<= 8'b00110100;
		7'b0100011: bcd_out<= 8'b00110101;
		7'b0100100: bcd_out<= 8'b00110110;
		7'b0100101: bcd_out<= 8'b00110111;
		7'b0100110: bcd_out<= 8'b00111000;
		7'b0100111: bcd_out<= 8'b00111001;
		7'b0101000: bcd_out<= 8'b01000000;
		7'b0101001: bcd_out<= 8'b01000001;
		7'b0101010: bcd_out<= 8'b01000010;
		7'b0101011: bcd_out<= 8'b01000011;
		7'b0101100: bcd_out<= 8'b01000100;
		7'b0101101: bcd_out<= 8'b01000101;
		7'b0101110: bcd_out<= 8'b01000110;
		7'b0101111: bcd_out<= 8'b01000111;
		7'b0110000: bcd_out<= 8'b01001000;
		7'b0110001: bcd_out<= 8'b01001001;
		7'b0110010: bcd_out<= 8'b01010000;
		7'b0110011: bcd_out<= 8'b01010001;
		7'b0110100: bcd_out<= 8'b01010010;
		7'b0110101: bcd_out<= 8'b01010011;
		7'b0110110: bcd_out<= 8'b01010100;
		7'b0110111: bcd_out<= 8'b01010101;
		7'b0111000: bcd_out<= 8'b01010110;
		7'b0111001: bcd_out<= 8'b01010111;
		7'b0111010: bcd_out<= 8'b01011000;
		7'b0111011: bcd_out<= 8'b01011001;
		7'b0111100: bcd_out<= 8'b01100000;
		7'b0111101: bcd_out<= 8'b01100001;
		7'b0111110: bcd_out<= 8'b01100010;
		7'b0111111: bcd_out<= 8'b01100011;
		7'b1000000: bcd_out<= 8'b01100100;
		7'b1000001: bcd_out<= 8'b01100101;
		7'b1000010: bcd_out<= 8'b01100110;
		7'b1000011: bcd_out<= 8'b01100111;
		7'b1000100: bcd_out<= 8'b01101000;
		7'b1000101: bcd_out<= 8'b01101001;
		7'b1000110: bcd_out<= 8'b01110000;
		7'b1000111: bcd_out<= 8'b01110001;
		7'b1001000: bcd_out<= 8'b01110010;
		7'b1001001: bcd_out<= 8'b01110011;
		7'b1001010: bcd_out<= 8'b01110100;
		7'b1001011: bcd_out<= 8'b01110101;
		7'b1001100: bcd_out<= 8'b01110110;
		7'b1001101: bcd_out<= 8'b01110111;
		7'b1001110: bcd_out<= 8'b01111000;
		7'b1001111: bcd_out<= 8'b01111001;
		7'b1010000: bcd_out<= 8'b10000000;
		7'b1010001: bcd_out<= 8'b10000001;
		7'b1010010: bcd_out<= 8'b10000010;
		7'b1010011: bcd_out<= 8'b10000011;
		7'b1010100: bcd_out<= 8'b10000100;
		7'b1010101: bcd_out<= 8'b10000101;
		7'b1010110: bcd_out<= 8'b10000110;
		7'b1010111: bcd_out<= 8'b10000111;
		7'b1011000: bcd_out<= 8'b10001000;
		7'b1011001: bcd_out<= 8'b10001001;
		7'b1011010: bcd_out<= 8'b10010000;
		7'b1011011: bcd_out<= 8'b10010001;
		7'b1011100: bcd_out<= 8'b10010010;
		7'b1011101: bcd_out<= 8'b10010011;
		7'b1011110: bcd_out<= 8'b10010100;
		7'b1011111: bcd_out<= 8'b10010101;
		7'b1100000: bcd_out<= 8'b10010110;
		7'b1100001: bcd_out<= 8'b10010111;
		7'b1100010: bcd_out<= 8'b10011000;
		7'b1100011: bcd_out<= 8'b10011001;
		default:
			bcd_out<= 8'b11101110;
	endcase
endmodule 