// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
// Created on Fri Jun 19 00:06:55 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module teste_fsm (
    input reset, input clock, input sign);

    enum int unsigned { state1=0, state2=1 } fstate, reg_fstate;

    always_ff @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always_comb begin
        if (reset) begin
            reg_fstate <= state1;
        end
        else begin
            case (fstate)
                state1: begin
                    if (sign)
                        reg_fstate <= state2;
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    if (sign)
                        reg_fstate <= state1;
                    else
                        reg_fstate <= state2;
                end
                default: begin
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // teste_fsm
